package VGA_config is

type VGA_config_t is record
  width  : natural; -- W: width
  height : natural; -- H: height
  rate   : natural; -- R: refresh rate
  clk    : natural; -- C: pixel clock (KHz)
  hpulse : natural; -- hS: horizontal sync pulse
  hfront : natural; -- hF: horizontal front porch
  hback  : natural; -- hB: horizontal back porch
  vpulse : natural; -- vS: vertical sync pulse
  vfront : natural; -- vF: vertical front porch
  vback  : natural; -- vB: vertical back porch
  hpol   : boolean; -- hP: inverted horizontal sync polarity?
  vpol   : boolean; -- hP: inverted vertical sync polarity?
end record;

--  PULSE FRONT LENGTH BACK
--   __                     __
-- _|  |XXXXXXX________XXXX|

type VGA_configs_t is array (natural range <>) of VGA_config_t;
constant VGA_configs : VGA_configs_t(0 to 61) := (
--           W      H     R        C    hS    hF    hB  vS    vF   vB      hP      vP
   0 => (  640,   350,   70,   25175,   96,   48,   16,  2,   60,  37,  false,   true ),
   1 => (  640,   350,   85,   31500,   64,   96,   32,  3,   60,  32,  false,   true ),
   2 => (  640,   400,   70,   25175,   96,   48,   16,  2,   35,  12,   true,  false ),
   3 => (  640,   400,   85,   31500,   64,   96,   32,  3,   41,   1,   true,  false ),
   4 => (  640,   480,   60,   25175,   96,   48,   16,  2,   33,  10,   true,   true ),
   5 => (  640,   480,   73,   31500,   40,  128,   24,  2,   29,   9,   true,   true ),
   6 => (  640,   480,   75,   31500,   64,  120,   16,  3,   16,   1,   true,   true ),
   7 => (  640,   480,   85,   36000,   56,   80,   56,  3,   25,   1,   true,   true ),
   8 => (  640,   480,  100,   43160,   64,  104,   40,  3,   25,   1,   true,  false ),
   9 => (  720,   400,   85,   35500,   72,  108,   36,  3,   42,   1,   true,  false ),
  10 => (  768,   576,   60,   34960,   80,  104,   24,  3,   17,   1,   true,  false ),
  11 => (  768,   576,   72,   42930,   80,  112,   32,  3,   21,   1,   true,  false ),
  12 => (  768,   576,   75,   45510,   80,  120,   40,  3,   22,   1,   true,  false ),
  13 => (  768,   576,   85,   51840,   80,  120,   40,  3,   25,   1,   true,  false ),
  14 => (  768,   576,  100,   62570,   80,  128,   48,  3,   31,   1,   true,  false ),
  15 => (  800,   600,   56,   36000,   72,  128,   24,  2,   22,   1,  false,  false ),
  16 => (  800,   600,   60,   40000,  128,   88,   40,  4,   23,   1,  false,  false ),
  17 => (  800,   600,   75,   49500,   80,  160,   16,  3,   21,   1,  false,  false ),
  18 => (  800,   600,   72,   50000,  120,   64,   56,  6,   23,  37,  false,  false ),
  19 => (  800,   600,   85,   56250,   64,  152,   32,  3,   27,   1,  false,  false ),
  20 => (  800,   600,  100,   68180,   88,  136,   48,  3,   32,   1,   true,  false ),
  21 => ( 1024,   768,   43,   44900,  176,   56,    8,  8,   41,   0,  false,  false ),
  22 => ( 1024,   768,   60,   65000,  136,  160,   24,  6,   29,   3,   true,   true ),
  23 => ( 1024,   768,   70,   75000,  136,  144,   24,  6,   29,   3,   true,   true ),
  24 => ( 1024,   768,   75,   78800,   96,  176,   16,  3,   28,   1,  false,  false ),
  25 => ( 1024,   768,   85,   94500,   96,  208,   48,  3,   36,   1,  false,  false ),
  26 => ( 1024,   768,  100,  113310,  112,  184,   72,  3,   42,   1,   true,  false ),
  27 => ( 1152,   864,   75,  108000,  128,  256,   64,  3,   32,   1,  false,  false ),
  28 => ( 1152,   864,   85,  119650,  128,  200,   72,  3,   39,   1,   true,  false ),
  29 => ( 1152,   864,  100,  143470,  128,  208,   80,  3,   47,   1,   true,  false ),
  30 => ( 1152,   864,   60,   81620,  120,  184,   64,  3,   27,   1,   true,  false ),
  31 => ( 1280,  1024,   60,  108000,  112,  248,   48,  3,   38,   1,  false,  false ),
  32 => ( 1280,  1024,   75,  135000,  144,  248,   16,  3,   38,   1,  false,  false ),
  33 => ( 1280,  1024,   85,  157500,  160,  224,   64,  3,   44,   1,  false,  false ),
  34 => ( 1280,  1024,  100,  190960,  144,  240,   96,  3,   57,   1,   true,  false ),
  35 => ( 1280,   800,   60,   83460,  136,  200,   64,  3,   24,   1,   true,  false ),
  36 => ( 1280,   960,   60,  102100,  136,  216,   80,  3,   30,   1,   true,  false ),
  37 => ( 1280,   960,   72,  124540,  136,  224,   88,  3,   37,   1,   true,  false ),
  38 => ( 1280,   960,   75,  129860,  136,  224,   88,  3,   38,   1,   true,  false ),
  39 => ( 1280,   960,   85,  148500,  160,  224,   64,  3,   47,   1,  false,  false ),
  40 => ( 1280,   960,  100,  178990,  144,  240,   96,  3,   53,   1,   true,  false ),
  41 => ( 1368,   768,   60,   85860,  144,  216,   72,  3,   23,   1,   true,  false ),
  42 => ( 1400,  1050,   60,  122610,  152,  240,   88,  3,   33,   1,   true,  false ),
  43 => ( 1400,  1050,   72,  149340,  152,  248,   96,  3,   40,   1,   true,  false ),
  44 => ( 1400,  1050,   75,  155850,  152,  248,   96,  3,   42,   1,   true,  false ),
  45 => ( 1400,  1050,   85,  179260,  152,  256,  104,  3,   49,   1,   true,  false ),
  46 => ( 1400,  1050,  100,  214390,  152,  264,  112,  3,   58,   1,   true,  false ),
  47 => ( 1440,   900,   60,  106470,  152,  232,   80,  3,   28,   1,   true,  false ),
  48 => ( 1600,  1200,   60,  162000,  192,  304,   64,  3,   46,   1,  false,  false ),
  49 => ( 1600,  1200,   65,  175500,  192,  304,   64,  3,   46,   1,  false,  false ),
  50 => ( 1600,  1200,   70,  189000,  192,  304,   64,  3,   46,   1,  false,  false ),
  51 => ( 1600,  1200,   75,  202500,  192,  304,   64,  3,   46,   1,  false,  false ),
  52 => ( 1600,  1200,   85,  229500,  192,  304,   64,  3,   46,   1,  false,  false ),
  53 => ( 1600,  1200,  100,  280640,  176,  304,  128,  3,   67,   1,   true,  false ),
  54 => ( 1680,  1050,   60,  147140,  184,  288,  104,  3,   33,   1,   true,  false ),
  55 => ( 1792,  1344,   60,  204800,  200,  328,  128,  3,   46,   1,   true,  false ),
  56 => ( 1792,  1344,   75,  261000,  216,  352,   96,  3,   69,   1,   true,  false ),
  57 => ( 1856,  1392,   60,  218300,  224,  352,   96,  3,   43,   1,   true,  false ),
  58 => ( 1856,  1392,   75,  288000,  224,  352,  128,  3,  104,   1,   true,  false ),
  59 => ( 1920,  1200,   60,  193160,  208,  336,  128,  3,   38,   1,   true,  false ),
  60 => ( 1920,  1440,   60,  234000,  208,  344,  128,  3,   56,   1,   true,  false ),
  61 => ( 1920,  1440,   75,  297000,  224,  352,  144,  3,   56,   1,   true,  false )
);

end VGA_config;
